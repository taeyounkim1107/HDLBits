module top_module(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);
	wire one, two;
    add16 inst1(a[15:0], b[15:0], 0, sum[15:0], one);
    add16 inst2(a[31:16], b[31:16], one, sum[31:16], two);
    
endmodule
